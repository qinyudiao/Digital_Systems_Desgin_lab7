`timescale 1ns / 10ps

module clockdiv(count_val, clk100Mhz, slowClk);
  input clk100Mhz; //fast clock
  input [27:0] count_val;
  output reg slowClk; //slow clock

  reg[27:0] counter;

  initial begin
    counter = 0;
    slowClk = 0;
  end

  always @ (posedge clk100Mhz)
  begin
    if(counter == count_val) begin
      counter <= 1;
      slowClk <= ~slowClk;
    end
    else begin
      counter <= counter + 1;
    end
  end

endmodule
